module Decoder_5to32(rd, rs1, rs2, Reg_rs1, Reg_rs2, en);  
input [4:0] rd, rs1, rs2; 
input en; 
output [31:0] Reg_rs1, Reg_rs2;
reg Reg_rs1, Reg_rs2; 
always @(rd or rs1 or rs2 or en)   begin 
if (en == 1'b1) 
case ( {rd,rs1,rs2} ) 
	5'b00000: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000000;
	5'b00001: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000001;
	5'b00010: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000010;
	5'b00011: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000011;
	5'b00100: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000100;
	5'b00101: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000101;
	5'b00110: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000110;
	5'b00111: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000000111;
	5'b01000: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001000;
	5'b01001: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001001;
	5'b01010: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001010;
	5'b01011: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001011;
	5'b01100: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001100;
	5'b01101: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001101;
	5'b01110: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001110;
	5'b01111: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000001111;
	5'b10000: {Reg_rs1, Reg_rs2} = 32'b00000000000000000000000000010000;
	default: {Reg_rs1, Reg_rs2} = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx; 
endcase 
if (en == 0) {Reg_rs1, Reg_rs2} = 32'b11111111111111111111111111111111; 
end 
endmodule